Test file for vhdl