Test file for vhd